module reciever_reader(offset_out, pwm_input, clk);
output offset_out;
input pwm_input;
input clk;

endmodule