module reciever_reader(offset_out, pwm_input);
output offset_out;
input pwm_input;

endmodule