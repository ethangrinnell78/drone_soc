module motor_offset_summer(motor_total_offset, pitch_offset, roll_offset, yaw_offset, throttle_offset, clk);
output motor_total_offset;
input pitch_offset;
input roll_offset;
input yaw_offset;
input throttle_offset;
input clk;

endmodule